`include "block_ram_pkg.sv"
`include "block_ram_if.sv"
