`ifndef AWIDTH
	`define AWIDTH 8
`endif 
`ifndef DWIDTH
	`define DWIDTH 8
`endif 
`ifndef MEM_DEPTH
	`define MEM_DEPTH 256
`endif 
